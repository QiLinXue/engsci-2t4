module hello_world ;

initial begin
  $display ("Hello World by Deepak");
   #10  $finish;
end

endmodule // End of Module hello_world